module top (
    output wifi_gpio0
);
    assign wifi_gpio0 = 1'b1;
endmodule
